** Profile: "Amp Diff-Time"  [ D:\PROJETPLURY\CARTE\Simulation\pp-amp diff-time.sim ] 

** Creating circuit file "pp-amp diff-time.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB ".\pp.lib" 
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.003 0 0.00003 
.STEP PARAM Gain LIST 10K, 20k 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\pp-Amp Diff.net" 


.END
